//gate level modelling
//and gate

//start module
module andGate(a,b,c);

//i/o ports
input a,b;
output c;

//intantiate primitive
and o (c,a,b);

//end module
endmodule
