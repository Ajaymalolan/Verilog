//gate level modelling
//not gate

//start module
module notGate(a,c);

//i/o ports
input a;
output c;

//intantiate primitive
not o (c,a);

//end module
endmodule
